`timescale 1ns/100ps
module tb_pe_conv_8x8();

reg clk = 0;
reg [127:0]in;
reg [17:0]filter;
wire [71:0]out;


always #5 clk=~clk;
top_pe_8x8 top_pe_8x80(clk,in,filter,out);

initial begin
	in[1:0]=1;in[3:2]=1;in[5:4]=0;in[7:6]=1;in[9:8]=1;in[11:10]=0;in[13:12]=0;in[15:14]=1;
	in[17:16]=0;in[19:18]=0;in[21:20]=1;in[23:22]=1;in[25:24]=1;in[27:26]=1;in[29:28]=1;in[31:30]=0;
	in[33:32]=1;in[35:34]=0;in[37:36]=0;in[39:38]=0;in[41:40]=1;in[43:42]=1;in[45:44]=0;in[47:46]=1;
	in[49:48]=0;in[51:50]=0;in[53:52]=0;in[55:54]=1;in[57:56]=0;in[59:58]=1;in[61:60]=0;in[63:62]=1;
	in[65:64]=1;in[67:66]=1;in[69:68]=0;in[71:70]=1;in[73:72]=0;in[75:74]=0;in[77:76]=1;in[79:78]=0;
	in[81:80]=0;in[83:82]=1;in[85:84]=1;in[87:86]=0;in[89:88]=1;in[91:90]=1;in[93:92]=0;in[95:94]=1;
	in[97:96]=1;in[99:98]=1;in[101:100]=1;in[103:102]=0;in[105:104]=1;in[107:106]=1;in[109:108]=0;in[111:110]=1;
	in[113:112]=1;in[115:114]=1;in[117:116]=0;in[119:118]=1;in[121:120]=0;in[123:122]=1;in[125:124]=1;in[127:126]=0;
	

	filter[1:0]=0;filter[3:2]=0;filter[5:4]=0;
	filter[7:6]=0;filter[9:8]=1;filter[11:10]=0;
	filter[13:12]=0;filter[15:14]=0;filter[17:16]=0;
	
	
	//$display("%d, %d, %d \n %d, %d, %d, \n %d, %d, %d",out[8:0],out[17:9],out[26:18],out[35:27],out[44:36],out[53:45],out[62:54],out[71:63],out[80:72]);
	
	
	
end
endmodule
